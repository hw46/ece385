module ripple_adder (
	input  logic  [7:0] a, 
    input  logic  [7:0] b,
	input  logic   m,
	input  logic   fn,//function select, add is 0, sub is 1
	
	output logic  [8:0] s,
	output logic   cout
);

	/* TODO
		*
		* Insert code here to implement a ripple adder.
		* Your code should be completly combinational (don't use always_ff or always_latch).
		* Feel free to create sub-modules or other files. */
	
logic c1,c2;
//logic [7:0] a_select; 
logic [7:0] b_select;
assign b_select = b ^ {8{fn}}; //invert B when fn = 1

		adder4 FA0 (.A (a[3:0]), .B (b_select[3:0]), .c_in(fn), .S (s[3:0]), .c_out (c1));
		adder4 FA1 (.A (a[7:4]), .B (b_select[7:4]), .c_in (c1), .S (s[7:4]), .c_out (c2));
		full_adder FA2 (.x (a[7]), .y (b_select[7]), .z (c2), .s (s[8]), .c (cout)); //calculate sign bit


endmodule



module full_adder (input x, y, z,
                   output s, c);
assign s = x^y^z;
assign c = (x&y)|(y&z)|(x&z);

endmodule


module adder4(input logic [3:0] A,B,
              input logic c_in,
              output logic [3:0]S,
              output logic c_out);
logic c1,c2,c3;
full_adder FA0 (.x (A[0]), .y (B[0]), .z (c_in), .s (S[0]), .c (c1));
full_adder FA1 (.x (A[1]), .y (B[1]), .z (c1), .s (S[1]), .c (c2));
full_adder FA2 (.x (A[2]), .y (B[2]), .z (c2), .s (S[2]), .c (c3));
full_adder FA3 (.x (A[3]), .y (B[3]), .z (c3), .s (S[3]), .c (c_out));              
              
endmodule

module ctrlx (input logic Clk,
              input logic load,
              input logic Reset,
              input logic in,
              output logic out);
 always_ff @(posedge Clk)
 begin
 if(Reset)out <= 1'b0;
 else out <= load ? in : out;
 end     
endmodule